module simd()
/*
make a mem file 
ALU can do only MAC, for 1 word of data, try to make this floating point
you can write another module to rearrange data
here, optimize things for matrix multiplication, do saturation and clipping calculations
*/

endmodule